LIBRARY ieee;
    USE ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    
    LIBRARY work;
    USE work.common.all;
    
    entity rom is
        port (address:  in  unsigned(7 downto 0);
              data_out: out bus_16_bit := (others => '1')
            );
    end entity rom;
    
    architecture behavior of rom is
    
    CONSTANT prom: bus_16_bit_vector(255 downto 0) := (
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1111111111111111",
"1010000000001010",
"1101101111001000",
"1100101100000000",
"0110101100010000",
"0110000100100000",
"1100000000000001",
"1010000010111101",
"0101000001000000",
"0101000100100000",
"1110001111000100",
"0110001110110000",
"0000001100001011",
"0001000100001011",
"0100010000000001",
"0100001000001010",
"0100000100001010",
"0100000000000000",
"1100000100000010",
"0100000100000000",
"1010000010111000",
"0110101100000000",
"0100000001100100",
"0100000100000001",
"1110000010110111",
"0110000010110000",
"0100000001100100",
"1100000100000100",
"1100000000000101",
"0000000100000001",
"0000000000000000",
"1010000010101110",
"0000101100001011",
"0001110000001011",
"0110110010110000",
"0100110000000000",
"0000000100000010",
"0000000000000010",
"1001101110101100",
"1110101110101100",
"0110101111000000",
"1010000010100011",
"0101101111000000",
"1101100010100010",
"0000110000010100",
"0001000100010100",
"0110000100000000",
"0100000100000000",
"1010000010011110",
"0001000000010100",
"1001001110011011",
"0000001100001010",
"1010000010010011",
"0110010001010000",
"0101000000110000",
"1001010010010111",
"0000010000001001",
"0100010100000001",
"0100001100001010",
"1010000010001100",
"0110010000110000",
"0101000000110000",
"1001010010010000",
"0100000000000000",
"0000010000001000",
"0100001100000001",
"0000101100010100",
"0001000100010100",
"0110000100000000",
"0100000100000000",
"1010000010001000",
"0001000000010100",
"1001001110000101",
"0000001100000111",
"1010000001111101",
"0110010001010000",
"0101000000110000",
"1001010010000001",
"0000010000000110",
"0100010100000001",
"0100001100001010",
"1010000001110110",
"0110010000110000",
"0101000000110000",
"1001010001111010",
"0100000000000000",
"0000010000000101",
"0100001100000001",
"1100000000000011",
"0000000000000100",
"1100000000000110",
"1100000000000111",
"0000000000000011",
"1010000000011111",
"1100000100000100",
"1100000000000101",
"0100000000000000",
"0100000100000001",
"0001110000000111",
"0001101100000110",
"0001101000000101",
"1010000001101010",
"0100000100000010",
"0001110000001010",
"0001101100001001",
"0001101000001000",
"1001110101100110",
"1100000100000010",
"1100000000000011",
"0000000100000010",
"0000000000000010",
"1010000001011110",
"0000000100000001",
"0000000000000000",
"1001110001011100",
"0111110000000000",
"0100000000000001",
"0100010000000000",
"0100001100000001",
"0101110001000000",
"1010000001010110",
"0100010000000001",
"0100001100000000",
"0101110000110000",
"1101011001010011",
"1100101100000001",
"0100101100000000",
"1010000001001101",
"1001000001001100",
"0110000010110000",
"0100000000001010",
"0100100000000001",
"0100011100000000",
"0101101101110000",
"1010000001001000",
"0100100000000000",
"0100011100000001",
"0101101110000000",
"1101010101000101",
"1100101000000000",
"0100101000000000",
"1010000000111111",
"1001000000111110",
"0110000010100000",
"0100000000001010",
"0100011000000001",
"0100010100000000",
"0101101001010000",
"1010000000111010",
"0100011000000000",
"0100010100000001",
"0101101001100000",
"1101010000110111",
"0100110100000000",
"0000110000000111",
"0000101100000110",
"0000101000000101",
"1010000000110010",
"0100110100000001",
"0000110000001010",
"0000101100001001",
"0000101000001000",
"1101011100101110",
"1100000100000110",
"1100000000000111",
"0000000100000010",
"0000000000000010",
"1010000000100110",
"0000000100000001",
"0000000000000000",
"1101100000100100",
"1101101101101110",
"0100010000000000",
"0100001100000001",
"0100100000000001",
"0100011100000000",
"1010000000011111",
"0100100000000000",
"0100011100000001",
"1101010100011011",
"0100011000000001",
"0100010100000000",
"1010000000010111",
"0100011000000000",
"0100010100000001",
"1101010000010101",
"0001000000001010",
"0001000000001001",
"0001000000001000",
"0001000000000111",
"0001000000000110",
"0001000000000101",
"0100000000000000",
"0001000000000100",
"0100000000001110",
"0001000000000011",
"0100000000001101",
"0001000000000010",
"0100000000001100",
"0001000000000001",
"0100000000001011",
"0001000000000000",
"0100000000001010"
);
    
    begin
    
    main: process(address)
    begin
        data_out <= prom(to_integer(address));
    end process main;
    
    end architecture behavior;